module ram(
	input clk,
	input ram_en,
	input ram_load,
    input stack_load,
    input mar_stack,
    input[11:0] mar,
    input[15:0] sp_out,
	input[15:0] bus,
	output[15:0] out
);

/*

0001MMMMMMMMMMMM	LDW
0010MMMMMMMMMMMM	STW
0011MMMMMMMMMMMM	ADD
0100MMMMMMMMMMMM	ADC
0101MMMMMMMMMMMM	SUB
0110MMMMMMMMMMMM	SBB
0111MMMMMMMMMMMM	MOD
1000MMMMMMMMMMMM	AND
1001MMMMMMMMMMMM	OR
1010MMMMMMMMMMMM	XOR
1011MMMMMMMMMMMM	JMP
1100MMMMMMMMMMMM	JPZ
1101MMMMMMMMMMMM	JPC
1110MMMMMMMMMMMM	JPS
1111MMMMMMMMMMMM	CAL
	
ZZZZ01SSSSSSSSSS	MSW
ZZZZ10SSSSSSSSSS	POP
ZZZZ11SSSSSSSSSS	RET
	
ZZZZZZ___001BBBB	BWS
ZZZZZZ___010BBBB	BWC
ZZZZZZ___011BBBB	BWJ
ZZZZZZ___100BBBB	BOS
ZZZZZZ___101BBBB	BOC
ZZZZZZ___110BBBB	BIJ
ZZZZZZ___111BBBB	BSL
	
ZZZZZZZZZZZZ0000	NOP
ZZZZZZZZZZZZ0001	INC
ZZZZZZZZZZZZ0010	DEC
ZZZZZZZZZZZZ0011	RTL
ZZZZZZZZZZZZ0100	RTR
ZZZZZZZZZZZZ0101	NOT
ZZZZZZZZZZZZ0110	COM
ZZZZZZZZZZZZ0111	LDP
ZZZZZZZZZZZZ1000	STP
ZZZZZZZZZZZZ1001	MWO
ZZZZZZZZZZZZ1010	MIW
ZZZZZZZZZZZZ1011	CLW
ZZZZZZZZZZZZ1100	CLO
ZZZZZZZZZZZZ1101	
ZZZZZZZZZZZZ1110	PSH
ZZZZZZZZZZZZ1111	RST

Z: unused opcode space
M: memory adress
S: distance above SP
B: bit in register

*/

reg[15:0] ram[0:12'b111111111111];

integer i;
initial begin
	$readmemb("program.bin", ram);
end

reg[15:0] out;
always @(posedge clk) begin
    if (ram_en) begin
		out <= ram[mar];
	end if (ram_load) begin
		ram[mar] <= bus;
    end if (stack_load) begin
        ram[sp_out] <= bus;
    end
end

endmodule